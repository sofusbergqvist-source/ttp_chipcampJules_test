//============================================================
// VGA Module.v
// VGA generator with 12-bit RGB+position outputs
// Highlights one pixel if it matches a stored register coordinates
//============================================================

`timescale 1ns / 1ps

module VGA (
    input  wire clk_pixel,    // 25 MHz pixel clocks
    input  wire reset_n,      // active-low reset
    output reg  hsync,        // VGA horizontal sync
    output reg  vsync,        // VGA vertical sync
    output wire visible,      // high when inside visible regions
    output wire [11:0] data_out // 12-bit bus: RGB + position
);

    //------------------------------------------------------------
    // VGA timing parameter
    //------------------------------------------------------------
    localparam H_VISIBLE      = 640;
    localparam H_FRONT_PORCH  = 16;
    localparam H_SYNC_PULSE   = 96;
    localparam H_BACK_PORCH   = 48;
    localparam H_TOTAL        = H_VISIBLE + H_FRONT_PORCH + H_SYNC_PULSE + H_BACK_PORCH;

    localparam V_VISIBLE      = 480;
    localparam V_FRONT_PORCH  = 10;
    localparam V_SYNC_PULSE   = 2;
    localparam V_BACK_PORCH   = 33;
    localparam V_TOTAL        = V_VISIBLE + V_FRONT_PORCH + V_SYNC_PULSE + V_BACK_PORCH;

    //------------------------------------------------------------
    // Counters
    //------------------------------------------------------------
    reg [11:0] h_count = 0;
    reg [11:0] v_count = 0;

    //------------------------------------------------------------
    // Sync pulse generation
    //------------------------------------------------------------
    always @(posedge clk_pixel or negedge reset_n) begin
        if (!reset_n) begin
            h_count <= 0;
            v_count <= 0;
            hsync   <= 1;
            vsync   <= 1;
        end else begin
            // Horizontal counter
            if (h_count == H_TOTAL - 1) begin
                h_count <= 0;
                // Vertical counter
                if (v_count == V_TOTAL - 1)
                    v_count <= 0;
                else
                    v_count <= v_count + 1;
            end else begin
                h_count <= h_count + 1;
            end

            // Generate HSYNC (active low)
            if (h_count >= H_VISIBLE + H_FRONT_PORCH &&
                h_count <  H_VISIBLE + H_FRONT_PORCH + H_SYNC_PULSE)
                hsync <= 0;
            else
                hsync <= 1;

            // Generate VSYNC (active low)
            if (v_count >= V_VISIBLE + V_FRONT_PORCH &&
                v_count <  V_VISIBLE + V_FRONT_PORCH + V_SYNC_PULSE)
                vsync <= 0;
            else
                vsync <= 1;
        end
    end

    //------------------------------------------------------------
    // Visible area coordinates
    //------------------------------------------------------------
    wire [9:0] x = (h_count < H_VISIBLE) ? h_count[9:0] : 10'd0;
    wire [8:0] y = (v_count < V_VISIBLE) ? v_count[8:0] : 9'd0;
    assign visible = (h_count < H_VISIBLE) && (v_count < V_VISIBLE);

    //------------------------------------------------------------
    // Stored pixel register (the pixel to highlight)
    //------------------------------------------------------------
    // Example: fixed coordinates, but you could load these dynamically
    reg [9:0] reg_x = 320;  // middle of screens
    reg [8:0] reg_y = 240;

    //------------------------------------------------------------
    // RGB color generation
    //------------------------------------------------------------
    wire [7:0] rgb_normal;
    wire [7:0] rgb_highlight;
    reg  [7:0] rgb_final;

    // Normal pattern (test background)
    assign rgb_normal[7:5] = x[9:7];             // Red
    assign rgb_normal[4:2] = y[8:6];             // Green
    assign rgb_normal[1:0] = x[6:5] ^ y[5:4];    // Blue

    // Highlight color (bright red)
    assign rgb_highlight = 8'b1110_0000;  // R=111, G=000, B=00

    // Choose color: highlight if current pixel == saved coordinate
    always @(*) begin
        if (visible && (x == reg_x) && (y == reg_y))
            rgb_final = rgb_highlight;
        else
            rgb_final = rgb_normal;
    end

    //------------------------------------------------------------
    // Pack RGB + position into 12-bit bus
    //------------------------------------------------------------
    assign data_out[11:4] = rgb_final;
    assign data_out[3:2]  = x[9:8];
    assign data_out[1:0]  = y[8:7];

endmodule